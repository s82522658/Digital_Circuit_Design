module BRICK(
	clk,
	col,
	row,
	b_col,
	b_row,
	brick
);
input clk;
input [10:0] col,row,b_col,b_row;
output brick;

wire [0:86*87-1] m_brick={
	87'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	87'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	87'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	87'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	87'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	87'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	87'b000000000000000000000000110000000000000000000000000000000000001000000000000000000000000,
	87'b000000000000000000000000111000000000000000000000000000000000011000000000000000000000000,
	87'b000000000000000000000000111100000000000000000000000000000000011000000000000000000000000,
	87'b000000000000000000000000111110000000000000000000000000000000111000000000000000000000000,
	87'b000000000000000000000000111111000000000000000000000000000001111000000000000000000000000,
	87'b000000000000000000000000111111110000000000000000000000000011111000000000000000000000000,
	87'b000000000000000000000000111111111000000000000000000000000111111000000000000000000000000,
	87'b000000000000000000000000111111111100000000000000000000011111111000000000000000000000000,
	87'b000000000000000000000000111111111110000000000000000000011111111100000000000000000000000,
	87'b000000000000000000000000111111111111100000000000000000111111111100000000000000000000000,
	87'b000000000000000000000001111111111111100000000000000001111111111100000000000000000000000,
	87'b000000000000000000000001111111111100000000000000000011111111111100000000000000000000000,
	87'b000000000000000000000001111111110000000000000000001111111111111100000000000000000000000,
	87'b000000000000000000000001111111100000001111111111001111111111111100000000000000000000000,
	87'b000000000000000000000001111110000011111111111111001111111111111100000000000000000000000,
	87'b000000000000000000000001111000011111111111111111101111111111111100000000000000000000000,
	87'b000000000000000000000001110000111111111111111111111111111111111100000000000000000000000,
	87'b000000000000000000000001100011111111111111111111111111111111111100000000000000000000000,
	87'b000000000000000000000000000111111111111111111111111111111111111100000000000000000000000,
	87'b000000000000000000000000001111111111111111111111111011111111111100000000000000000000000,
	87'b000000000000000000000000011111111111111111111111111110111111111000000000000000000000000,
	87'b000000000000000000000000111111111111111111111111111111101110000000000000000000000000000,
	87'b000000000000000000000001111111111111111111111111111111110000000000000000000000000000000,
	87'b000000000000000000000001111111111111111111111111111111111110001100000000000000000000000,
	87'b000000000000000000000011111111111111111111111111111111111111111110000000000000000000000,
	87'b000000000000000000000011111111111111111111111111111111111111111100000000000000000000000,
	87'b000000000000000000000111111111111111111111111111111111111111111001111000000000000000000,
	87'b000000000000000111000111111111111111111111111111111111111111111011111111100000000000000,
	87'b000000000011111111001111111111111111111111111111111111111111110111111111111110000000000,
	87'b000000001111111110001111111111111111111111111111111111111111111111111111111111111000000,
	87'b000000000111111110011111111111111111111111111111111111111111111111111111111111111110000,
	87'b000000000011111110011111111111111100111111001111111111111111111111111111111111111100000,
	87'b000000000001111110011111111111111100111111001111111111111111111111111111111111111000000,
	87'b000000000000111100011111111111111111111111101111111111111111011111111111111111100000000,
	87'b000000000000011100111111111111111111111111111111111111111111011111111111111111000000000,
	87'b000000000000001100111111111111111111111111111111111111111111011111111111111110000000000,
	87'b000000000000001000111111111111111111111111111111111111111111101111111111111100000000000,
	87'b000000000000000000111111111111111111111111111111111111111111101111111111111000000000000,
	87'b000000000000000000111111111111111111111111111111111111111111110111111111110000000000000,
	87'b000000000000000000111111111111111111111111111111111111111111110011111111100000000000000,
	87'b000000000000000000111111111111111111111111111111111111111111111000111111000000000000000,
	87'b000000000000000000111111111111111111111111111111111111111111111100000000000000000000000,
	87'b000000000000000000111111111111111111111111111111111111111111111110000000000000000000000,
	87'b000000000000000000111111111111111111111111111111111111111111111111110000000000000000000,
	87'b000000000000000000011111111111111111111111111111111111111111111111111000000000000000000,
	87'b000000000000000000011111111111111111111111111111111111111111111111111000000000000000000,
	87'b000000000000000000011111111111111111111111111111111111111111111111110000000000000000000,
	87'b000000000000000000001111111111111111111111111111111111111111111111110000000000000000000,
	87'b000000000000000000001111111111111111111111111111111111111111111111100000000000000000000,
	87'b000000000000000000000111111111111111111111111111111111111111111111100000000000000000000,
	87'b000000000000000000000111111111111111111111111111111111111111111111100000000000000000000,
	87'b000000000000000000000011111111111111111111111111111111111111111111111000000000000000000,
	87'b000000000000000000000011111111111111111111111111111111111111111111111110000000000000000,
	87'b000000000000000000000001111111111111111111111111111111111111111111111110000000000000000,
	87'b000000000000000000000000111111111111111111111111111111111111111111111111000000000000000,
	87'b000000000000000000000000011111111111111111111111111111111111111111111111100000000000000,
	87'b000000000000000000000000111111111111111111111111111111111111111111111111110000000000000,
	87'b000000000000000000000000111111111111111111111111111111111111111111111111110000000000000,
	87'b000000000000000000000001111111111111111111111111111111111111111111111111110000000000000,
	87'b000000000000000000000001111111111111111111111111111111111111111111111111100000000000000,
	87'b000000000000000000000001111111111111111111111111111111111111111111111111111000000000000,
	87'b000000000000000000000001111111111111111111111111111111111111111111111111111000000000000,
	87'b000000000000000000000011111111111111111111111111111111111111111111111111111000000000000,
	87'b000000000000000000000011111111111111111111111111111111111111111111111111100000000000000,
	87'b000000000000000000000011111111111111111111111111111111111111111111111111100000000000000,
	87'b000000000000000000000011111111111111111111111111111111111111111111111111111000000000000,
	87'b000000000000000000000011111111111111111111111111111111111111111111111111100000000000000,
	87'b000000000000000000000011111111111111111111111111111111111111111111111111111000000000000,
	87'b000000000000000000000011111111111111111111111111111111111111111111111111111000000000000,
	87'b000000000000000000000001111111111111111111111111111111111111111111111111111000000000000,
	87'b000000000000000000000001111111111111111111111111111111111111111111111111110000000000000,
	87'b000000000000000000000001111111111111111111111111111111111111111111111111100000000000000,
	87'b000000000000000000000000111111111111111111111111111111111111111111111111000000000000000,
	87'b000000000000000000000000011111111111111111111111111111111111111111111111000000000000000,
	87'b000000000000000000000000011111111111111111111111111111111111111111111100000000000000000,
	87'b000000000000000000000000001111111111111111111111111111111111111111110000000000000000000,
	87'b000000000000000000000000000111111111111111111111111111111111111111100000000000000000000,
	87'b000000000000000000000000000000111111111111111111111111111111111110000000000000000000000,
	87'b000000000000000000000000000000001111111111111111111111111111111000000000000000000000000,
	87'b000000000000000000000000000000000000000111111111111111111100000000000000000000000000000
};
assign brick = (m_brick[(row-b_row)*87+(col-b_col)])? 1:0;
/*
//brick
always@(posedge clk) begin
	if((row-b_row)>=37 & (row-b_row)<=39 & (col-b_col)>=34 & (col-b_col)<=43 & !m_brick[(row-b_row)*87+(col-b_col)])brick<=3'b000;//eyes black
	else if(m_brick[(row-b_row)*87+(col-b_col)]) brick<=3'b010;//body green
	else brick<=3'b000;//black
end
*/
endmodule