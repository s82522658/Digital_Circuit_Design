`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:02:53 12/28/2015 
// Design Name: 
// Module Name:    Bricker 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////


module GAMEOVER(clk,col,row,gg
    );
input clk;
input [10:0]col,row;
output reg [2:0]gg;
reg [49:0]line1,line2,line3,line4,line5,line6,line7,line8,line9,line10,line11,line12,line13,line14,line15,line16,line17,line18,line19,line20
,line21,line22,line23,line24,line25,line26,line27,line28,line29,line30,line31,line32,line33,line34,line35,line36,line37,line38,line39,line40,line41;
reg [9:0] col_e;
reg flag;

always@(*)begin
	if(col > 140 & col <=190) col_e = 190; 
	else if(col > 200 & col <=250) col_e = 250;
	else if(col > 260 & col <=310) col_e = 310;
	else if(col > 320 & col <=370) col_e = 370;
	else if(col > 430 & col <=480) col_e = 480;
	else if(col > 490 & col <=540) col_e = 540;
	else if(col > 550 & col <=600) col_e = 600;
	else if(col > 610 & col <=660) col_e = 660;
	else col_e = 0;
end



always@(*)begin
	case (col_e)
		190:begin 
			line1  = 50'b00000000000000000111111111111111111000000000000000;
			line2  = 50'b00000000000001111111111111111111111111111100000000;
			line3  = 50'b00000000001111111111111111111111111111111111000000;
			line4  = 50'b00000000111111111111111111111111111111111111000000;
			line5  = 50'b00000011111111111111111000000001111111111111000000;
			line6  = 50'b00000111111111111111000000000000001111111111000000;
			line7  = 50'b00001111111111111110000000000000000111111111000000;
			line8  = 50'b00011111111111111100000000000000000011111111000000;
			line9  = 50'b00011111111111111000000000000000000011111111000000;
			line10 = 50'b00111111111111110000000000000000000001111111000000;
			line11 = 50'b00111111111111100000000000000000000001111111000000;
			line12 = 50'b01111111111111000000000000000000000001111111000000;
			line13 = 50'b01111111111111000000000000000000000001111111000000;
			line14 = 50'b01111111111111000000000000000000000000000000000000;
			line15 = 50'b11111111111111000000000000000000000000000000000000;
			line16 = 50'b11111111111110000000000000000000000000000000000000;
			line17 = 50'b11111111111110000000000000000000000000000000000000;
			line18 = 50'b11111111111110000000000000000000000000000000000000;
			line19 = 50'b11111111111110000000000000000000000000000000000000;
			line20 = 50'b11111111111110000000000000000000000000000000000000;
			line21 = 50'b11111111111110000000000000000000000000000000000000;
			line22 = 50'b11111111111110000000000001111111111111111111111111;
			line23 = 50'b11111111111110000000000001111111111111111111111111;
			line24 = 50'b11111111111110000000000001111111111111111111111111;
			line25 = 50'b11111111111110000000000001111111111111111111111111;
			line26 = 50'b11111111111110000000000000000001111111111111111100;
			line27 = 50'b11111111111110000000000000000000011111111111110000;
			line28 = 50'b01111111111111000000000000000000011111111111100000;
			line29 = 50'b01111111111111000000000000000000011111111111100000;
			line30 = 50'b01111111111111000000000000000000011111111111100000;
			line31 = 50'b00111111111111100000000000000000011111111111100000;
			line32 = 50'b00111111111111100000000000000000011111111111100000;
			line33 = 50'b00011111111111110000000000000000011111111111100000;
			line34 = 50'b00011111111111111000000000000000011111111111100000;
			line35 = 50'b00001111111111111100000000000000011111111111100000;
			line36 = 50'b00000111111111111111000000000001111111111111100000;
			line37 = 50'b00000011111111111111111100011111111111111111100000;
			line38 = 50'b00000000111111111111111111111111111111111111100000;
			line39 = 50'b00000000011111111111111111111111111111111111100000;
			line40 = 50'b00000000000011111111111111111111111100000000000000;
			line41 = 50'b00000000000000000111111111111110000000000000000000;
		end
		250:begin 
			line1  = 50'b00000000000000000000000000000000000000000000000000;
			line2  = 50'b00000000000000000001111111111110000000000000000000;
			line3  = 50'b00000000000000000001111111111111000000000000000000;
			line4  = 50'b00000000000000000011111111111111000000000000000000;
			line5  = 50'b00000000000000000011111111111111100000000000000000;
			line6  = 50'b00000000000000000111111111111111100000000000000000;
			line7  = 50'b00000000000000000111111111111111100000000000000000;
			line8  = 50'b00000000000000001111111111111111110000000000000000;
			line9  = 50'b00000000000000001111111111111111110000000000000000;
			line10 = 50'b00000000000000001111111111111111111000000000000000;
			line11 = 50'b00000000000000011111111111111111111000000000000000;
			line12 = 50'b00000000000000011111111111111111111000000000000000;
			line13 = 50'b00000000000000011111111111111111111100000000000000;
			line14 = 50'b00000000000000111111111111111111111100000000000000;
			line15 = 50'b00000000000000111111111111111111111110000000000000;
			line16 = 50'b00000000000001111111111111111111111110000000000000;
			line17 = 50'b00000000000001111111111100111111111111000000000000;
			line18 = 50'b00000000000011111111111100111111111111000000000000;
			line19 = 50'b00000000000011111111111100111111111111100000000000;
			line20 = 50'b00000000000011111111111100011111111111100000000000;
			line21 = 50'b00000000000111111111111000011111111111100000000000;
			line22 = 50'b00000000000111111111111000001111111111110000000000;
			line23 = 50'b00000000001111111111110000001111111111110000000000;
			line24 = 50'b00000000001111111111110000001111111111110000000000;
			line25 = 50'b00000000001111111111110000000111111111111000000000;
			line26 = 50'b00000000011111111111100000000111111111111000000000;
			line27 = 50'b00000000011111111111111111111111111111111100000000;
			line28 = 50'b00000000111111111111111111111111111111111100000000;
			line29 = 50'b00000000111111111111111111111111111111111100000000;
			line30 = 50'b00000000111111111111111111111111111111111110000000;
			line31 = 50'b00000001111111111111111111111111111111111110000000;
			line32 = 50'b00000001111111111111111111111111111111111111000000;
			line33 = 50'b00000011111111111111111111111111111111111111000000;
			line34 = 50'b00000011111111111111111111111111111111111111100000;
			line35 = 50'b00000111111111111100000000000000111111111111100000;
			line36 = 50'b00000111111111111100000000000000111111111111100000;
			line37 = 50'b00000111111111111000000000000000011111111111110000;
			line38 = 50'b00001111111111111000000000000000011111111111110000;
			line39 = 50'b00001111111111111000000000000000001111111111111000;
			line40 = 50'b00011111111111110000000000000000001111111111111000;
			line41 = 50'b00000000000000000000000000000000000000000000000000;
		end
		310:begin 
			line1  = 50'b00000000000000000000000000000000000000000000000000;
			line2  = 50'b11111111111110000000000000000000000001111111111111;
			line3  = 50'b11111111111110000000000000000000000001111111111111;
			line4  = 50'b00001111111111000000000000000000000011111111111100;
			line5  = 50'b00000111111111100000000000000000000011111111110000;
			line6  = 50'b00000111111111100000000000000000000111111111100000;
			line7  = 50'b00000011111111110000000000000000000111111111100000;
			line8  = 50'b00000011111111110000000000000000001111111111100000;
			line9  = 50'b00000011111111110000000000000000001111111111100000;
			line10 = 50'b00000011111111111000000000000000001111111111100000;
			line11 = 50'b00000011111111111000000000000000011111111111100000;
			line12 = 50'b00000011111111111000000000000000011110111111100000;
			line13 = 50'b00000011111111111100000000000000111110111111100000;
			line14 = 50'b00000011111111111100000000000000111100111111100000;
			line15 = 50'b00000011110111111110000000000001111100111111100000;
			line16 = 50'b00000011110111111110000000000001111000111111100000;
			line17 = 50'b00000011110011111111000000000001111000111111100000;
			line18 = 50'b00000011110011111111000000000011110000111111100000;
			line19 = 50'b00000011110001111111100000000011110000111111100000;
			line20 = 50'b00000011110001111111100000000111110000111111100000;
			line21 = 50'b00000011110000111111110000000111100000111111100000;
			line22 = 50'b00000011110000111111110000001111100000111111100000;
			line23 = 50'b00000011110000011111111000001111000000111111100000;
			line24 = 50'b00000011110000011111111000011111000000111111100000;
			line25 = 50'b00000011110000001111111100011110000000111111100000;
			line26 = 50'b00000011110000001111111100111110000000111111100000;
			line27 = 50'b00000011110000000111111110111110000000111111100000;
			line28 = 50'b00000011110000000111111110111100000000111111100000;
			line29 = 50'b00000011110000000011111111111100000000111111100000;
			line30 = 50'b00000011110000000011111111111000000000111111100000;
			line31 = 50'b00000011110000000001111111111000000000111111100000;
			line32 = 50'b00000011110000000001111111110000000000111111100000;
			line33 = 50'b00000011110000000001111111110000000000111111100000;
			line34 = 50'b00000011110000000000111111110000000000111111100000;
			line35 = 50'b00000011110000000000111111100000000000111111100000;
			line36 = 50'b00000111110000000000011111000000000000111111100000;
			line37 = 50'b00001111111000000000011111000000000001111111110000;
			line38 = 50'b01111111111111000000001110000000001111111111111110;
			line39 = 50'b11111111111111100000001110000000011111111111111111;
			line40 = 50'b11111111111111100000000100000000011111111111111111;
			line41 = 50'b00000000000000000000000000000000000000000000000000;
		end
		370:begin 
			line1  = 50'b00000000111111111111111111111111111111111000000000;
			line2  = 50'b00000000111111111111111111111111111111111000000000;
			line3  = 50'b00000000111111111111111111111111111111111000000000;
			line4  = 50'b00000000000011111111111111111111111111111000000000;
			line5  = 50'b00000000000001111111000000000000000111111000000000;
			line6  = 50'b00000000000001111111000000000000000011111000000000;
			line7  = 50'b00000000000001111111000000000000000001111000000000;
			line8  = 50'b00000000000001111111000000000000000001111000000000;
			line9  = 50'b00000000000001111111000000000000000000111000000000;
			line10 = 50'b00000000000001111111000000000000000000111000000000;
			line11 = 50'b00000000000001111111000000000000000000000000000000;
			line12 = 50'b00000000000001111111000000000000000000000000000000;
			line13 = 50'b00000000000001111111000000000000000110000000000000;
			line14 = 50'b00000000000001111111000000000000001110000000000000;
			line15 = 50'b00000000000001111111000000000000001110000000000000;
			line16 = 50'b00000000000001111111000000000000001110000000000000;
			line17 = 50'b00000000000001111111000000000000011110000000000000;
			line18 = 50'b00000000000001111111000000000000011110000000000000;
			line19 = 50'b00000000000001111111111111111111111110000000000000;
			line20 = 50'b00000000000001111111111111111111111110000000000000;
			line21 = 50'b00000000000001111111111111111111111110000000000000;
			line22 = 50'b00000000000001111111111111111111111110000000000000;
			line23 = 50'b00000000000001111111000000000000011110000000000000;
			line24 = 50'b00000000000001111111000000000000001110000000000000;
			line25 = 50'b00000000000001111111000000000000001110000000000000;
			line26 = 50'b00000000000001111111000000000000001110000000000000;
			line27 = 50'b00000000000001111111000000000000000110000000000000;
			line28 = 50'b00000000000001111111000000000000000000000000000000;
			line29 = 50'b00000000000001111111000000000000000000000000000000;
			line30 = 50'b00000000000001111111000000000000000000000111000000;
			line31 = 50'b00000000000001111111000000000000000000001111000000;
			line32 = 50'b00000000000001111111000000000000000000001110000000;
			line33 = 50'b00000000000001111111000000000000000000011110000000;
			line34 = 50'b00000000000001111111000000000000000000011110000000;
			line35 = 50'b00000000000001111111000000000000000000111110000000;
			line36 = 50'b00000000000001111111000000000000000001111100000000;
			line37 = 50'b00000000000001111111000000000000001111111100000000;
			line38 = 50'b00000000000011111111111111111111111111111100000000;
			line39 = 50'b00000000111111111111111111111111111111111100000000;
			line40 = 50'b00000000111111111111111111111111111111111000000000;
			line41 = 50'b00000000111111111111111111111111111111111000000000;
		end
		480:begin 
			line1  = 50'b00000000000000000000000000000000000000000000000000;
			line2  = 50'b00000000000000000000111111111111000000000000000000;
			line3  = 50'b00000000000000001111111111111111110000000000000000;
			line4  = 50'b00000000000000111111100000000111111100000000000000;
			line5  = 50'b00000000000011111110000000000000111111100000000000;
			line6  = 50'b00000000000111111100000000000000111111100000000000;
			line7  = 50'b00000000001111111000000000000000011111110000000000;
			line8  = 50'b00000000011111110000000000000000001111111000000000;
			line9  = 50'b00000000111111100000000000000000000111111100000000;
			line10 = 50'b00000000111111100000000000000000000011111110000000;
			line11 = 50'b00000001111111000000000000000000000011111110000000;
			line12 = 50'b00000001111111000000000000000000000011111111000000;
			line13 = 50'b00000011111111000000000000000000000001111111000000;
			line14 = 50'b00000011111111000000000000000000000001111111000000;
			line15 = 50'b00000011111111000000000000000000000001111111100000;
			line16 = 50'b00000111111110000000000000000000000001111111100000;
			line17 = 50'b00000111111110000000000000000000000001111111100000;
			line18 = 50'b00000111111110000000000000000000000001111111100000;
			line19 = 50'b00000111111110000000000000000000000001111111100000;
			line20 = 50'b00000111111110000000000000000000000001111111100000;
			line21 = 50'b00000111111110000000000000000000000001111111100000;
			line22 = 50'b00000111111110000000000000000000000001111111100000;
			line23 = 50'b00000111111110000000000000000000000001111111100000;
			line24 = 50'b00000111111110000000000000000000000001111111100000;
			line25 = 50'b00000111111110000000000000000000000001111111100000;
			line26 = 50'b00000111111110000000000000000000000001111111100000;
			line27 = 50'b00000111111111000000000000000000000001111111100000;
			line28 = 50'b00000011111111000000000000000000000001111111000000;
			line29 = 50'b00000011111111000000000000000000000011111110000000;
			line30 = 50'b00000011111111000000000000000000000011111110000000;
			line31 = 50'b00000001111111100000000000000000000011111110000000;
			line32 = 50'b00000001111111100000000000000000000111111100000000;
			line33 = 50'b00000000111111110000000000000000000111111100000000;
			line34 = 50'b00000000111111110000000000000000001111111000000000;
			line35 = 50'b00000000001111111000000000000000011111110000000000;
			line36 = 50'b00000000000111111100000000000000111111100000000000;
			line37 = 50'b00000000000011111111000000000001111111000000000000;
			line38 = 50'b00000000000000111111100000000011111110000000000000;
			line39 = 50'b00000000000000001111111111111111110000000000000000;
			line40 = 50'b00000000000000000001111111111111000000000000000000;
			line41 = 50'b00000000000000000000000000000000000000000000000000;
		end
		540:begin 
			line1  = 50'b00111111111111111111111000000000011111111111111000;
			line2  = 50'b00111111111111111111111000000000011111111111111000;
			line3  = 50'b00111111111111111111111000000000011111111111111000;
			line4  = 50'b00000111111111111111000000000000000011111111100000;
			line5  = 50'b00000011111111111110000000000000000001111110000000;
			line6  = 50'b00000001111111111110000000000000000001111100000000;
			line7  = 50'b00000000111111111110000000000000000001111100000000;
			line8  = 50'b00000000111111111110000000000000000001111000000000;
			line9  = 50'b00000000011111111111000000000000000001111000000000;
			line10 = 50'b00000000011111111111000000000000000011110000000000;
			line11 = 50'b00000000001111111111100000000000000011110000000000;
			line12 = 50'b00000000001111111111100000000000000111100000000000;
			line13 = 50'b00000000001111111111110000000000000111100000000000;
			line14 = 50'b00000000000111111111110000000000001111000000000000;
			line15 = 50'b00000000000111111111110000000000001111000000000000;
			line16 = 50'b00000000000011111111111000000000001111000000000000;
			line17 = 50'b00000000000011111111111000000000011110000000000000;
			line18 = 50'b00000000000001111111111100000000011110000000000000;
			line19 = 50'b00000000000001111111111100000000111100000000000000;
			line20 = 50'b00000000000000111111111110000000111100000000000000;
			line21 = 50'b00000000000000111111111110000000111100000000000000;
			line22 = 50'b00000000000000111111111111000001111000000000000000;
			line23 = 50'b00000000000000011111111111000001111000000000000000;
			line24 = 50'b00000000000000011111111111000011110000000000000000;
			line25 = 50'b00000000000000001111111111100011110000000000000000;
			line26 = 50'b00000000000000001111111111100111100000000000000000;
			line27 = 50'b00000000000000000111111111110111100000000000000000;
			line28 = 50'b00000000000000000111111111110111100000000000000000;
			line29 = 50'b00000000000000000011111111111111000000000000000000;
			line30 = 50'b00000000000000000011111111111111000000000000000000;
			line31 = 50'b00000000000000000011111111111110000000000000000000;
			line32 = 50'b00000000000000000001111111111110000000000000000000;
			line33 = 50'b00000000000000000001111111111100000000000000000000;
			line34 = 50'b00000000000000000000111111111100000000000000000000;
			line35 = 50'b00000000000000000000111111111100000000000000000000;
			line36 = 50'b00000000000000000000011111111000000000000000000000;
			line37 = 50'b00000000000000000000011111111000000000000000000000;
			line38 = 50'b00000000000000000000001111110000000000000000000000;
			line39 = 50'b00000000000000000000001111110000000000000000000000;
			line40 = 50'b00000000000000000000000111100000000000000000000000;
			line41 = 50'b00000000000000000000000111100000000000000000000000;
		end
		600:begin 
			line1  = 50'b00000000111111111111111111111111111111111000000000;
			line2  = 50'b00000000111111111111111111111111111111111000000000;
			line3  = 50'b00000000111111111111111111111111111111111000000000;
			line4  = 50'b00000000000011111111111111111111111111111000000000;
			line5  = 50'b00000000000001111111000000000000000111111000000000;
			line6  = 50'b00000000000001111111000000000000000011111000000000;
			line7  = 50'b00000000000001111111000000000000000001111000000000;
			line8  = 50'b00000000000001111111000000000000000001111000000000;
			line9  = 50'b00000000000001111111000000000000000000111000000000;
			line10 = 50'b00000000000001111111000000000000000000111000000000;
			line11 = 50'b00000000000001111111000000000000000000000000000000;
			line12 = 50'b00000000000001111111000000000000000000000000000000;
			line13 = 50'b00000000000001111111000000000000000110000000000000;
			line14 = 50'b00000000000001111111000000000000001110000000000000;
			line15 = 50'b00000000000001111111000000000000001110000000000000;
			line16 = 50'b00000000000001111111000000000000001110000000000000;
			line17 = 50'b00000000000001111111000000000000011110000000000000;
			line18 = 50'b00000000000001111111000000000000011110000000000000;
			line19 = 50'b00000000000001111111111111111111111110000000000000;
			line20 = 50'b00000000000001111111111111111111111110000000000000;
			line21 = 50'b00000000000001111111111111111111111110000000000000;
			line22 = 50'b00000000000001111111111111111111111110000000000000;
			line23 = 50'b00000000000001111111000000000000011110000000000000;
			line24 = 50'b00000000000001111111000000000000001110000000000000;
			line25 = 50'b00000000000001111111000000000000001110000000000000;
			line26 = 50'b00000000000001111111000000000000001110000000000000;
			line27 = 50'b00000000000001111111000000000000000110000000000000;
			line28 = 50'b00000000000001111111000000000000000000000000000000;
			line29 = 50'b00000000000001111111000000000000000000000000000000;
			line30 = 50'b00000000000001111111000000000000000000000111000000;
			line31 = 50'b00000000000001111111000000000000000000001111000000;
			line32 = 50'b00000000000001111111000000000000000000001110000000;
			line33 = 50'b00000000000001111111000000000000000000011110000000;
			line34 = 50'b00000000000001111111000000000000000000011110000000;
			line35 = 50'b00000000000001111111000000000000000000111110000000;
			line36 = 50'b00000000000001111111000000000000000001111100000000;
			line37 = 50'b00000000000001111111000000000000001111111100000000;
			line38 = 50'b00000000000011111111111111111111111111111100000000;
			line39 = 50'b00000000111111111111111111111111111111111100000000;
			line40 = 50'b00000000111111111111111111111111111111111000000000;
			line41 = 50'b00000000111111111111111111111111111111111000000000;
		end
		660:begin 
			line1  = 50'b00000000000000000000000000000000000000000000000000;
			line2  = 50'b01111111111111111111111111111111100000000000000000;
			line3  = 50'b01111111111111111111111111111111111110000000000000;
			line4  = 50'b01111111111111111111111111111111111111100000000000;
			line5  = 50'b01111111111111111111111111111111111111110000000000;
			line6  = 50'b01111111111111111111111111111111111111111000000000;
			line7  = 50'b00000001111111111110000000111111111111111000000000;
			line8  = 50'b00000001111111111110000000001111111111111100000000;
			line9  = 50'b00000001111111111110000000000111111111111100000000;
			line10 = 50'b00000001111111111110000000000111111111111100000000;
			line11 = 50'b00000001111111111110000000000111111111111100000000;
			line12 = 50'b00000001111111111110000000000111111111111100000000;
			line13 = 50'b00000001111111111110000000000111111111111100000000;
			line14 = 50'b00000001111111111110000000000111111111111100000000;
			line15 = 50'b00000001111111111110000000001111111111111000000000;
			line16 = 50'b00000001111111111110000000001111111111111000000000;
			line17 = 50'b00000001111111111110000000111111111111110000000000;
			line18 = 50'b00000001111111111110000011111111111111100000000000;
			line19 = 50'b00000001111111111111111111111111111111000000000000;
			line20 = 50'b00000001111111111111111111111111111000000000000000;
			line21 = 50'b00000001111111111111111111111110000000000000000000;
			line22 = 50'b00000001111111111111111111111111000000000000000000;
			line23 = 50'b00000001111111111111111111111111100000000000000000;
			line24 = 50'b00000001111111111111111111111111110000000000000000;
			line25 = 50'b00000001111111111110111111111111111000000000000000;
			line26 = 50'b00000001111111111110011111111111111100000000000000;
			line27 = 50'b00000001111111111110001111111111111110000000000000;
			line28 = 50'b00000001111111111110000111111111111110000000000000;
			line29 = 50'b00000001111111111110000111111111111111000000000000;
			line30 = 50'b00000001111111111110000011111111111111100000000000;
			line31 = 50'b00000001111111111110000001111111111111110000000000;
			line32 = 50'b00000001111111111110000000111111111111111000000000;
			line33 = 50'b00000001111111111110000000011111111111111100000000;
			line34 = 50'b00000001111111111110000000001111111111111100000000;
			line35 = 50'b00000001111111111110000000000111111111111111000000;
			line36 = 50'b00000111111111111111100000000111111111111111110000;
			line37 = 50'b01111111111111111111111110000011111111111111111110;
			line38 = 50'b01111111111111111111111110000001111111111111111110;
			line39 = 50'b01111111111111111111111110000001111111111111111110;
			line40 = 50'b01111111111111111111111110000000111111111111111110;
			line41 = 50'b00000000000000000000000000000000000000000000000000;
		end
		default:begin
			line1  = 0;
			line2  = 0;
			line3  = 0;
			line4  = 0;
			line5  = 0;
			line6  = 0;
			line7  = 0;
			line8  = 0;
			line9  = 0;
			line10 = 0;
			line11 = 0;
			line12 = 0;
			line13 = 0;
			line14 = 0;
			line15 = 0;
			line16 = 0;
			line17 = 0;
			line18 = 0;
			line19 = 0;
			line20 = 0;
			line21 = 0;
			line22 = 0;
			line23 = 0;
			line24 = 0;
			line25 = 0;
			line26 = 0;
			line27 = 0;
			line28 = 0;
			line29 = 0;
			line30 = 0;
			line31 = 0;
			line32 = 0;
			line33 = 0;
			line34 = 0;
			line35 = 0;
			line36 = 0;
			line37 = 0;
			line38 = 0;
			line39 = 0;
			line40 = 0;
			line41 = 0;		
		end
	endcase
end


always@(*)begin
	if(row >=280 & row <= 320 & ~(col_e==0) )begin
		case(row)
			280 : flag = line1  [col_e-col];
			281 : flag = line2  [col_e-col];
			282 : flag = line3  [col_e-col];
			283 : flag = line4  [col_e-col];
			284 : flag = line5  [col_e-col];
			285 : flag = line6  [col_e-col];
			286 : flag = line7  [col_e-col];
			287 : flag = line8  [col_e-col];
			288 : flag = line9  [col_e-col];
			289 : flag = line10 [col_e-col];
			290 : flag = line11 [col_e-col];
			291 : flag = line12 [col_e-col];
			292 : flag = line13 [col_e-col];
			293 : flag = line14 [col_e-col];
			294 : flag = line15 [col_e-col];
			295 : flag = line16 [col_e-col];
			296 : flag = line17 [col_e-col];
			297 : flag = line18 [col_e-col];
			298 : flag = line19 [col_e-col];
			299 : flag = line20 [col_e-col];
			300 : flag = line21 [col_e-col];
			301 : flag = line22 [col_e-col];
			302 : flag = line23 [col_e-col];
			303 : flag = line24 [col_e-col];
			304 : flag = line25 [col_e-col];
			305 : flag = line26 [col_e-col];
			306 : flag = line27 [col_e-col];
			307 : flag = line28 [col_e-col];
			308 : flag = line29 [col_e-col];
			309 : flag = line30 [col_e-col];
			310 : flag = line31 [col_e-col];
			311 : flag = line32 [col_e-col];
			312 : flag = line33 [col_e-col];
			313 : flag = line34 [col_e-col];
			314 : flag = line35 [col_e-col];
			315 : flag = line36 [col_e-col];
			316 : flag = line37 [col_e-col];
			317 : flag = line38 [col_e-col];
			318 : flag = line39 [col_e-col];
			319 : flag = line40 [col_e-col];
			320 : flag = line41 [col_e-col];
			default: flag = 0;
		endcase
	end
	else flag = 0;
end

always@(posedge clk)begin
	if(flag) gg <= 3'b100;
	else gg <= 3'b000;
end
	
endmodule 