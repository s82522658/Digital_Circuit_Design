module CANDY(
	clk,
	row,
	col,
	c_row,
	c_col,
	candy
);
input clk;
input [10:0] col,row,c_col,c_row;
//output reg [2:0] candy;
output   candy;
reg flag;
wire [0:80*84-1] m_candy ={
	84'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
	84'b1111111111111111111111111111111111111111111111111111111111111111111100000111111111111,
	84'b1111111111101111111111111111111111111111111111111111111111111111110000000001111111111,
	84'b1111111100000001111111111111111111111111111111111111111111111111100000000000011111111,
	84'b1111111000000000011111111111111110000000000000000111111111111111000000000000011111111,
	84'b1111110000000000001111111111110000000000000000000000011111111110000000000000001111111,
	84'b1111100000000000000111111110000000000000000000000000000111111100000000000000001111111,
	84'b1111000000000000000011111000000000000000000000000000000001111000000000000000001111111,
	84'b1111000000000000000001100000000000000000000000000000000000010000000000000000001111111,
	84'b1111000000000000000000000000000000000000000000000000000000000000000000000000001111111,
	84'b1111000000000000000000000000000000000000000000000000000000000000000000000000001111111,
	84'b1111000000000000000000000000000000000000000000000000000000000000000000000000001111111,
	84'b1111000000000000000000000000000000000000000000000000000000000000000000000000001111111,
	84'b1111000000000000000000000000000000000000000000000000000000000000000000000000011111111,
	84'b1111000000000000000000000000000000000000000000000000000000000000000000000000011111111,
	84'b1111100000000000000000000000000000000000000000000000000000000000000000000000111111111,
	84'b1111100000000000000000000000000000000000000000000000000000000000000000000000111111111,
	84'b1111110000000000000000000000000000000000000000000000000000000000000000000001111111111,
	84'b1111110000000000000000000000000000000000000000000000000000000000000000000001111111111,
	84'b1111111000000000000000000000000000000000000000000000000000000000000000000011111111111,
	84'b1111111100000000000000000000000000000000000000000000000000000000000000000011111111111,
	84'b1111111100000000000000000000000000000000000000000000000000000000000000000011111111111,
	84'b1111111110000000000000000000000000000000000000000000000000000000000000000001111111111,
	84'b1111111100000000000000000000000000000000000000000000000000000000000000000000111111111,
	84'b1111111000000000000000000000000000000000000000000000000000000000000000000000011111111,
	84'b1111111000000000000000111111000000000000000000000000001111110000000000000000011111111,
	84'b1111110000000000000000000000000000000011111110000000000000000000000000000000001111111,
	84'b1111110000000000000000000000000000001111111111000000000000000000000000000000001111111,
	84'b1111100000000000000000000000000000001111111111000000000000000000000000000000000111111,
	84'b1111100000000000000000000000000000001111111111000000000000000000000000000000000111111,
	84'b1111100000000000000000000000000000000111111111000000000000000000000000000000000011111,
	84'b1111000000000000000000000000000000000011111000000000000000000000000000000000000011111,
	84'b1111000000000000000000000000000000000000010000000000000000000000000000000000000011111,
	84'b1111000000000000000000000000000000000000010000000000000000000000000000000000000001111,
	84'b1111000000000000000000000000000000000000010000000000000000000000000000000000000001111,
	84'b1110000000000000000000000000000001000000110000001000000000000000000000000000000001111,
	84'b1110000000000000000000000000000001100000111000001000000000000000000000000000000001111,
	84'b1110000000000000000000000000000000111111111111110000000000000000000000000000000001111,
	84'b1110000000000000000000000000000000001111111111100000000000000000000000000000000001111,
	84'b1110000000000000000000000000000000001111111111100000000000000000000000000000000001111,
	84'b1110000000000000000000000000000000001111111111100000000000000000000000000000000001111,
	84'b1110000000000000000000000000000000001111111111000000000000000000000000000000000001111,
	84'b1110000000000000000000000000000000000111111111000000000000000000000000000000000001111,
	84'b1110000000000000000000000000000000000111111111000000000000000000000000000000000001111,
	84'b1110000000000000000000000000000000000111111111000000000000000000000000000000000001111,
	84'b1110000000000000000000000000000000000011111110000000000000000000000000000000000001111,
	84'b1110000000000000000000000000000000000001111100000000000000000000000000000000000001111,
	84'b1111000000000000000000000000000000000000000000000000000000000000000000000000000011111,
	84'b1111000000000000000000000000000000000000000000000000000000000000000000000000000011111,
	84'b1111000000000000000000000000000000000000000000000000000000000000000000000000000011111,
	84'b1111000000000000000000000000000000000000000000000000000000000000000000000000000011111,
	84'b1111100000000000000000000000000000000000000000000000000000000000000000000000000111111,
	84'b1111100000000000000000000000000000000000000000000000000000000000000000000000000111111,
	84'b1111100000000000000000000000000000000000000000000000000000000000000000000000001111111,
	84'b1111110000000000000000000000000000000000000000000000000000000000000000000000001111111,
	84'b1111110000000000000000000000000000000000000000000000000000000000000000000000011111111,
	84'b1111111000000000000000000000000000000000000000000000000000000000000000000000011111111,
	84'b1111111100000000000000000000000000000000000000000000000000000000000000000000111111111,
	84'b1111111100000000000000000000000000000000000000000000000000000000000000000000111111111,
	84'b1111111110000000000000000000000000000000000000000000000000000000000000000001111111111,
	84'b1111111111000000000000000000000000000000000000000000000000000000000000000011111111111,
	84'b1111111111000000000000000000000000000000000000000000000000000000000000000011111111111,
	84'b1111111111100000000000000000000000000000000000000000000000000000000000000111111111111,
	84'b1111111111110000000000000000000000000000000000000000000000000000000000001111111111111,
	84'b1111111111111000000000000000000000000000000000000000000000000000000000011111111111111,
	84'b1111111111111100000000000000000000000000000000000000000000000000000000111111111111111,
	84'b1111111111111110000000000000000000000000000000000000000000000000000001111111111111111,
	84'b1111111111111111000000000000000000000000000000000000000000000000000011111111111111111,
	84'b1111111111111111110000000000000000000000000000000000000000000000000111111111111111111,
	84'b1111111111111111111000000000000000000000000000000000000000000000001111111111111111111,
	84'b1111111111111111111110000000000000000000000000000000000000000000111111111111111111111,
	84'b1111111111111111111111000000000000000000000000000000000000000011111111111111111111111,
	84'b1111111111111111111111111000000000000000000000000000000000000111111111111111111111111,
	84'b1111111111111111111111111110000000000000000000000000000000111111111111111111111111111,
	84'b1111111111111111111111111111110000000000000000000000000111111111111111111111111111111,
	84'b1111111111111111111111111111111111000000000000000000111111111111111111111111111111111,
	84'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
	84'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
	84'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
	84'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111
};

assign candy = (!m_candy[(row-c_row)*84+(col-c_col)])? 1:0;//�給1 五��
/*
//candy
always@(posedge clk) begin
	if(!m_candy[(row-c_row)*84+(col-c_col)]) candy<=3'b101;//face pink
	else if((row-c_row)>=25 & (row-c_row)<=46 & (col-c_col)>=22 & (col-c_col)<=59 & flag) candy<=3'b100;//五� red
	else candy<= 3'b110;//ground yellow ?? 
end
*/
endmodule