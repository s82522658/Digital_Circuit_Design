`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:52:34 01/06/2017 
// Design Name: 
// Module Name:    RUNNING 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module running(
	clk,
	rst,
	VGA_RED,
	VGA_GREEN,
	VGA_BLUE,
	VGA_HSYNC,
	VGA_VSYNC,
    kclk,
    kdata,
	LCD_E,
	LCD_RS,
	LCD_RW,
	LCD_D,
    start_button
);

input clk,rst,kclk,kdata,start_button;
output VGA_RED,VGA_GREEN,VGA_BLUE,VGA_HSYNC,VGA_VSYNC;
output LCD_E,LCD_RS,LCD_RW;
output [3:0] LCD_D;
reg [103:0] row_a,row_b;
	

wire visible;
wire [10:0] col,row;
wire [2:0] bird;//bird enable
wire [1:0] tree;//tree enable
wire [2:0] back;//back color
wire  brick,brick1,brick2,brick3,brick4;//brick enable
wire candy;//candy enable
wire [90:0] gg_0,gg_1,gg_2,gg_3,gg_4,gg_5,gg_6,gg_7,gg_8,gg_9,gg_10,gg_11,gg_12,gg_13,gg_14,gg_15,gg_16,gg_17,gg_18,gg_19,gg_20,gg_21,gg_22,gg_23,gg_24,gg_25,gg_26,gg_27,gg_28,gg_29,gg_30,gg_31,gg_32,gg_33,gg_34,gg_35,gg_36,gg_37,gg_38,gg_39,gg_40,gg_41,gg_42,gg_43,gg_44,gg_45,gg_46,gg_47,gg_48,gg_49,gg_50,gg_51,gg_52,gg_53,gg_54,gg_55,gg_56,gg_57,gg_58,gg_59,gg_60,gg_61,gg_62,gg_63,gg_64,gg_65,gg_66,gg_67,gg_68,gg_69,gg_70,gg_71,gg_72,gg_73,gg_74,gg_75,gg_76,gg_77,gg_78,gg_79,gg_80,gg_81,gg_82,gg_83,gg_84,gg_85,gg_86,gg_87;
wire [115:0] g1,g2,g3,g4,g5,g6,g7,g8,g9,g10,g11,g12,g13,g14,g15,g16,g17,g18,g19,g20,g21,g22,g23,g24,g25,g26,g27,g28,g29,g30,g31,g32,g33,g34,g35,g36,g37,g38,g39,g40,g41,g42,g43,g44,g45,g46,g47,g48,g49,g50,g51,g52;
wire rele;
wire [10:0] c_row= 270;
wire check;
wire moon;
wire [2:0]gg,win;
wire rfd,rfd1;
wire [3:0]fractional,fractional1;
wire[7:0] quo,quo1;


reg c_state,n_state;
reg day;
reg [3:0] key_counter;
reg [21:0] key_reg;
reg [7:0] key_data;
reg [10:0] yb_cnt;
reg [1:0] yb_flag;
reg up_cho;
reg [2:0] color;
reg [10:0] pixel_col,pixel_row;
reg [10:0] bk_col,bk_col1,bk_col2,bk_col3,bk_col4,c_col;
reg [10:0] s_col,m_col;
reg [10:0] up_col;
reg [25:0] counter,cnt;
reg [5:0] random;
reg [4:0] bk_cho;
reg [5:0] bk_num;
reg [2:0] timer;
reg choose,choose2,choose3;
reg nnflag,nflag;
reg [10:0]gg_row;
integer gg_col = 120,g_col = 120,g_row = 449;
reg [1:0] move;// 0:rst 1:up 2:down
reg start,Flag;
reg [1:0]fg;
reg [26:0] halfseccnt;
reg halfsec;
reg gflag,gameover;
reg [2:0] life;
reg [3:0] t_invincible;
reg invincible;
reg c_cho;
reg blink;


parameter H_fp=919;
parameter H_bp=104;
parameter H_pw=1039;
parameter H_disp=904;
parameter V_fp=659;
parameter V_bp=23;
parameter V_pw=665;
parameter V_disp=623;
parameter SUN=0;
parameter MOON=1;

assign VGA_RED = color[2];
assign VGA_GREEN = color[1];
assign VGA_BLUE = color[0];
assign VGA_HSYNC=~(pixel_col >= H_fp & pixel_col < H_pw);
assign VGA_VSYNC=~(pixel_row >= V_fp & pixel_row < V_pw);
assign visible=( pixel_col>=H_bp & pixel_col<H_disp & pixel_row>=V_bp & pixel_row<V_disp );//timing of display 
assign col=pixel_col - H_bp;
assign row=pixel_row - V_bp;
/*
BRICK BR (
    .clk(clk), 
    .col(col), 
    .row(row), 
    .b_col(bk_col), 
    .b_row(414), //414~499
    .brick(brick)
    );	
BRICK B1 (
    .clk(clk), 
    .col(col), 
    .row(row), 
    .b_col(bk_col1), 
    .b_row(414), //414~499
    .brick(brick1)
    );	
BRICK B2 (
    .clk(clk), 
    .col(col), 
    .row(row), 
    .b_col(bk_col2), 
    .b_row(414), //414~499
    .brick(brick2)
    );	
BRICK B3 (
    .clk(clk), 
    .col(col), 
    .row(row), 
    .b_col(bk_col3), 
    .b_row(414), //414~499
    .brick(brick3)
    );	
BRICK B4 (
    .clk(clk), 
    .col(col), 
    .row(row), 
    .b_col(bk_col4), 
    .b_row(414), //414~499
    .brick(brick4)
    );
	*/

LCD L1 (
	.LCD_E(LCD_E),
    .LCD_RS(LCD_RS), 
    .LCD_RW(LCD_RW), 
    .LCD_D(LCD_D), 
	.row_a(row_a), 
	.clk(clk),
    .btn_s(rst)
    );		
CANDY c1 (
    .clk(clk), 
    .col(col), 
    .row(row), 
	.c_row(c_row), 
	.c_col(c_col),
    .candy(candy)
    );	
GAMEOVER instance_name (
    .clk(clk), 
    .col(col), 
    .row(row), 
    .gg(gg)
    );
	
WIN instance_name1 (
    .clk(clk), 
    .col(col), 
    .row(row), 
    .win(win)
    );
	
divi pass(
	.clk(clk), // input clk
	.rfd(rfd), // output rfd
	.dividend(bk_num), // input [15 : 0] dividend
	.divisor(10), // input [15 : 0] divisor
	.quotient(quo), // output [15 : 0] quotient
	.fractional(fractional)
	); 
divi remain(
	.clk(clk), // input clk
	.rfd(rfd1), // output rfd
	.dividend(20-bk_bum), // input [15 : 0] dividend
	.divisor(10), // input [15 : 0] divisor
	.quotient(quo1), // output [15 : 0] quotient
	.fractional(fractional1)
	);

/////////////////

//////board/////
//n_state,c_state
always@(posedge clk)begin
	c_state <= n_state;
	n_state <= kclk;
end
//key_reg
always@(posedge clk)begin
	case({c_state,n_state})
		2'b10 : begin 
			key_reg <= {kdata,key_reg[21:1]};
			if(key_counter >=10) key_counter <= 0;
			else key_counter <= key_counter +1;
		end
		default : key_reg <= key_reg;
	endcase
end

assign check = key_reg[1]^key_reg[2]^key_reg[3]^key_reg[4]^key_reg[5]^key_reg[6]^key_reg[7]^key_reg[8]^key_reg[9];
//yb_flag,start
always@(posedge clk or posedge rst)begin
	if(rst) begin yb_flag <= 2; start<=0; end
	else if( key_counter==0 && check == 1 )begin
		if( key_reg[8:1] == 8'hF0 ) yb_flag <= 2;
		else if(key_reg[19:12]==8'h75 ) yb_flag <= 0;
		else if(key_reg[19:12]==8'h72 ) yb_flag <= 1;
        else if(key_reg[19:12]==8'h5A ) start<=1;
		else begin yb_flag <= yb_flag; start<=start; end
	end
	else begin yb_flag <= yb_flag; start<=start; end
end


//-------halfsec------
always@ (posedge clk or posedge rst) begin
	halfseccnt<=(rst)?0:(halfseccnt<185000)?halfseccnt+1:0;
	halfsec<=(rst)?0:(halfseccnt==0)?~halfsec:halfsec;
end
//---------------------

///////nn/////////

assign gg_0 = 91'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign gg_1 = 91'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign gg_2 = 91'b0000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000;
assign gg_3 = 91'b0000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000;
assign gg_4 = 91'b0000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000;
assign gg_5 = 91'b0000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000;
assign gg_6 = 91'b0000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000;
assign gg_7 = 91'b0000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000;
assign gg_8 = 91'b0000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000;
assign gg_9 = 91'b0000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000;
assign gg_10 = 91'b0000000000000000000000000000000000000001111111111111111111111111110000000000000000000000000;
assign gg_11 = 91'b0000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000;
assign gg_12 = 91'b0000000000000000000000000000000000000111111111111111111111111111111100000000000000000000000;
assign gg_13 = 91'b0000000000000000000000000000000000000111111111111111111111111111111100000000000000000000000;
assign gg_14 = 91'b0000000000000000000000000000000000000111111111001111111110011111111110000000000000000000000;
assign gg_15 = 91'b0000000000000000000000000000000000000111111111001111111110011111111110000000000000000000000;
assign gg_16 = 91'b0000000000000000000000000000000000001111111110000111111100001111111110000000000000000000000;
assign gg_17 = 91'b0000000000000000000000000000000000001111111110000111111100001111111110000000000000000000000;
assign gg_18 = 91'b0000000000000000000000000000000000001111111111001111111110011111111111000000000000000000000;
assign gg_19 = 91'b0000000000000000000000000000000000001111111111001111111110011111111111000000000000000000000;
assign gg_20 = 91'b0000000000000000000000000000000000001111111111111111111111111111111111000000000000000000000;
assign gg_21 = 91'b0000000000000000000000000000000000001111111111111111111111111111111111000000000000000000000;
assign gg_22 = 91'b0000000000000000000000000000000000001111111111111111111111111111111110000000000000000000000;
assign gg_23 = 91'b0000000000000000000000000000000000001111111111111111111111111111111110000000000000000000000;
assign gg_24 = 91'b0000000000000000000000000000000000001111111111111111111111111111111110000000000000000000000;
assign gg_25 = 91'b0000000000000000000000000000000000001111111111111111111111111111111110000000000000000000000;
assign gg_26 = 91'b0000000000000000000000000000000000000111111111111111111111111111111100000000000000000000000;
assign gg_27 = 91'b0000000000000000000000000000000000000111111111111111111111111111111100000000000000000000000;
assign gg_28 = 91'b0000000000000000000000000001111100000011111111111111111111111111111100001111110000000000000;
assign gg_29 = 91'b0000000000000000000000000001111100000011111111111111111111111111111100001111110000000000000;
assign gg_30 = 91'b0000000000000000000000001111111111111001111111111111111111111111111111111111111110000000000;
assign gg_31 = 91'b0000000000000000000000001111111111111001111111111111111111111111111111111111111110000000000;
assign gg_32 = 91'b0000000000000000000000111111111111111111111111111100000000111111111111111111111111100000000;
assign gg_33 = 91'b0000000000000000000000111111111111111111111111111100000000111111111111111111111111100000000;
assign gg_34 = 91'b0000000000000000000001111111111111111111111111111000000000011111111111111111111111110000000;
assign gg_35 = 91'b0000000000000000000001111111111111111111111111111000000000011111111111111111111111110000000;
assign gg_36 = 91'b0000000000000000000001111111111111111111111111111100000000111111111110001111111111110000000;
assign gg_37 = 91'b0000000000000000000001111111111111111111111111111111111111111111111100011111111111110000000;
assign gg_38 = 91'b0000000000000000000001111111111111111111111111111111111111111111111110001111111111111000000;
assign gg_39 = 91'b0000000000000000000001111111111111000111111111111111111111111111111110011111111111111000000;
assign gg_40 = 91'b0000000000000000000001111111111110000111111111111100000000111111111111111111111111110000000;
assign gg_41 = 91'b0000000000000000000001111111111111000111111111111000000000011111111111111111111111110000000;
assign gg_42 = 91'b0000000000000000000001111111111111001111111111111000000000011111111111111111111111110000000;
assign gg_43 = 91'b0000000000000000000001111111111111111111111111111100000000111111111111111111111111110000000;
assign gg_44 = 91'b0000000000000000000000011111111111111111111111111111111111111111111111111111111111100000000;
assign gg_45 = 91'b0000000000000000000000011111111111111111111111111111111111111111111111111111111111100000000;
assign gg_46 = 91'b0000000000000000000000000111111111111111111111111111111111111111111111111111111110000000000;
assign gg_47 = 91'b0000000000000000000000000111111111111111111111111111111111111111111111111111111110000000000;
assign gg_48 = 91'b0000000000000000000000000000011111111111111111111111111111111111111111111111000000000000000;
assign gg_49 = 91'b0000000000000000000000000000011111111111111111111111111111111111111111111111000000000000000;
assign gg_50 = 91'b0000000000000000000000000000000000111111111111111111111111111111111111110000000000000000000;
assign gg_51 = 91'b0000000000000000000000000000000000111111111111111111111111111111111111110000000000000000000;
assign gg_52 = 91'b0000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000;
assign gg_53 = 91'b0000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000;
assign gg_54 = 91'b0000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000;
assign gg_55 = 91'b0000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000;
assign gg_56 = 91'b0000000000000000000000000000000000000001111111111111111111111111111000000000000000000000000;
assign gg_57 = 91'b0000000000000000000000000000000000000001111111111111111111111111111000000000000000000000000;
assign gg_58 = 91'b0000000000000000000000000000000000000111111111111111111111111111111100000000000000000000000;
assign gg_59 = 91'b0000000000000000000000000000000000000111111111111111111111111111111100000000000000000000000;
assign gg_60 = 91'b0000000000000000000000000000000000011111111111111111111111111111111111000000000000000000000;
assign gg_61 = 91'b0000000000000000000000000000000000011111111111111111111111111111111111000000000000000000000;
assign gg_62 = 91'b0000000000000000000000000000000000111111111111111111111111111111111111110000000000000000000;
assign gg_63 = 91'b0000000000000000000000000000000000111111111111111111111111111111111111110000000000000000000;
assign gg_64 = 91'b0000000000000000000000000000000011111111111111111111111111111111111111111000000000000000000;
assign gg_65 = 91'b0000000000000000000000000000000011111111111111111111111111111111111111111000000000000000000;
assign gg_66 = 91'b0000000000000000000000000000001111111111111111111111111111111111111111111110000000000000000;
assign gg_67 = 91'b0000000000000000000000000000001111111111111111111111111111111111111111111110000000000000000;
assign gg_68 = 91'b0000000000000000000000000000011111111111111111111111111111111111111111111111100000000000000;
assign gg_69 = 91'b0000000000000000000000000000011111111111111111111111111111111111111111111111100000000000000;
assign gg_70 = 91'b0000000000000000000000000001111111111111111111111111011111111111111111111111110000000000000;
assign gg_71 = 91'b0000000000000000000000000001111111111111111111111111011111111111111111111111110000000000000;
assign gg_72 = 91'b0000000000000000000000000011111111111111111111111110001111111111111111111111111000000000000;
assign gg_73 = 91'b0000000000000000000000000011111111111111111111111110001111111111111111111111111000000000000;
assign gg_74 = 91'b0000000000000000000000000011111111111111111111111000000011111111111111111111111000000000000;
assign gg_75 = 91'b0000000000000000000000000011111111111111111111111000000011111111111111111111111000000000000;
assign gg_76 = 91'b0000000000000000000000000011111111111111111111100000000000111111111111111111111000000000000;
assign gg_77 = 91'b0000000000000000000000000011111111111111111111100000000000111111111111111111111000000000000;
assign gg_78 = 91'b0000000000000000000000000011111111111111111110000000000000011111111111111111111000000000000;
assign gg_79 = 91'b0000000000000000000000000011111111111111111110000000000000011111111111111111111000000000000;
assign gg_80 = 91'b0000000000000000000000000011111111111111111100000000000000000111111111111111111000000000000;
assign gg_81 = 91'b0000000000000000000000000011111111111111111100000000000000000111111111111111111000000000000;
assign gg_82 = 91'b0000000000000000000000000000111111111111110000000000000000000001111111111111100000000000000;
assign gg_83 = 91'b0000000000000000000000000000111111111111110000000000000000000001111111111111100000000000000;
assign gg_84 = 91'b0000000000000000000000000000001111111111000000000000000000000000011111111110000000000000000;
assign gg_85 = 91'b0000000000000000000000000000001111111111000000000000000000000000011111111110000000000000000;
assign gg_86 = 91'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign gg_87 = 91'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//nnflag
always @(posedge clk) begin
	if(col > gg_col && col <= gg_col+91 && row > gg_row && row <=gg_row + 87)begin
		case(row-gg_row)
		0 : nnflag <= gg_0[col];
		1 : nnflag <= gg_1[col];
		2 : nnflag <= gg_2[col];
		3 : nnflag <= gg_3[col];
		4 : nnflag <= gg_4[col];
		5 : nnflag <= gg_5[col];
		6 : nnflag <= gg_6[col];
		7 : nnflag <= gg_7[col];
		8 : nnflag <= gg_8[col];
		9 : nnflag <= gg_9[col];
		10 : nnflag <= gg_10[col];
		11 : nnflag <= gg_11[col];
		12 : nnflag <= gg_12[col];
		13 : nnflag <= gg_13[col];
		14 : nnflag <= gg_14[col];
		15 : nnflag <= gg_15[col];
		16 : nnflag <= gg_16[col];
		17 : nnflag <= gg_17[col];
		18 : nnflag <= gg_18[col];
		19 : nnflag <= gg_19[col];
		20 : nnflag <= gg_20[col];
		21 : nnflag <= gg_21[col];
		22 : nnflag <= gg_22[col];
		23 : nnflag <= gg_23[col];
		24 : nnflag <= gg_24[col];
		25 : nnflag <= gg_25[col];
		26 : nnflag <= gg_26[col];
		27 : nnflag <= gg_27[col];
		28 : nnflag <= gg_28[col];
		29 : nnflag <= gg_29[col];
		30 : nnflag <= gg_30[col];
		31 : nnflag <= gg_31[col];
		32 : nnflag <= gg_32[col];
		33 : nnflag <= gg_33[col];
		34 : nnflag <= gg_34[col];
		35 : nnflag <= gg_35[col];
		36 : nnflag <= gg_36[col];
		37 : nnflag <= gg_37[col];
		38 : nnflag <= gg_38[col];
		39 : nnflag <= gg_39[col];
		40 : nnflag <= gg_40[col];
		41 : nnflag <= gg_41[col];
		42 : nnflag <= gg_42[col];
		43 : nnflag <= gg_43[col];
		44 : nnflag <= gg_44[col];
		45 : nnflag <= gg_45[col];
		46 : nnflag <= gg_46[col];
		47 : nnflag <= gg_47[col];
		48 : nnflag <= gg_48[col];
		49 : nnflag <= gg_49[col];
		50 : nnflag <= gg_50[col];
		51 : nnflag <= gg_51[col];
		52 : nnflag <= gg_52[col];
		53 : nnflag <= gg_53[col];
		54 : nnflag <= gg_54[col];
		55 : nnflag <= gg_55[col];
		56 : nnflag <= gg_56[col];
		57 : nnflag <= gg_57[col];
		58 : nnflag <= gg_58[col];
		59 : nnflag <= gg_59[col];
		60 : nnflag <= gg_60[col];
		61 : nnflag <= gg_61[col];
		62 : nnflag <= gg_62[col];
		63 : nnflag <= gg_63[col];
		64 : nnflag <= gg_64[col];
		65 : nnflag <= gg_65[col];
		66 : nnflag <= gg_66[col];
		67 : nnflag <= gg_67[col];
		68 : nnflag <= gg_68[col];
		69 : nnflag <= gg_69[col];
		70 : nnflag <= gg_70[col];
		71 : nnflag <= gg_71[col];
		72 : nnflag <= gg_72[col];
		73 : nnflag <= gg_73[col];
		74 : nnflag <= gg_74[col];
		75 : nnflag <= gg_75[col];
		76 : nnflag <= gg_76[col];
		77 : nnflag <= gg_77[col];
		78 : nnflag <= gg_78[col];
		79 : nnflag <= gg_79[col];
		80 : nnflag <= gg_80[col];
		81 : nnflag <= gg_81[col];
		82 : nnflag <= gg_82[col];
		83 : nnflag <= gg_83[col];
		84 : nnflag <= gg_84[col];
		85 : nnflag <= gg_85[col];
		86 : nnflag <= gg_86[col];
		87 : nnflag <= gg_87[col];
		endcase
	end
end

//---------�Ʀ檺����H---------
assign g1 = 116'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign g2 = 116'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign g3 = 116'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign g4 = 116'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign g5 = 116'b00000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000;
assign g6 = 116'b00000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000;
assign g7 = 116'b00000000000000000000000000000000000000111111111111111111111000000000000000000000000000000000000000000000000000000000;
assign g8 = 116'b00000000000000000000000000000000000011111111111111111111111100000000000000000000000000000000000000000000000000000000;
assign g9 = 116'b00000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000000000000000000000000;
assign g10 = 116'b00000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000000000000000000000000000;
assign g11 = 116'b00000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000;
assign g12 = 116'b00000000000000000000000000000000111111111111111110000111111111111100000000000000000000000000000000000000000000000000;
assign g13 = 116'b00000000000000000000000000000001111111111111111100000011111111111100000000000000000000000000000000000000000000000000;
assign g14 = 116'b00000000000000000000000000000011111111111111111100000011111111111110000000000000000000000000000000000000000000000000;
assign g15 = 116'b00000000000000000000000000000011111111111111111100000011111111111110000000000000000000000000000000000000000000000000;
assign g16 = 116'b00000000000000000000000000000111111111111111111100000111111111111111000000000000000000000000000000000000000000000000;
assign g17 = 116'b00000000000000000000000000000111111111111111111111001111111111111111000000000000000000000000000000000000000000000000;
assign g18 = 116'b00000000000000000000000000001111111111111111111111111111111111111111100000000000000000000000000000000000000000000000;
assign g19 = 116'b00000000000000000000000000001111111111111111111111111111111000011111100000000000000000000000000000000000000000000000;
assign g20 = 116'b00000000000000000000000000001111111111111111111111111111110011111111100000000000000000000000000000000000000000000000;
assign g21 = 116'b00000000000000000000000000001111111111111111111111111111100111001111100000000000000000000000000000000000000000000000;
assign g22 = 116'b00000000000000000000000000011111111111111111111111111111101111001111100000000000000000000000000000000000000000000000;
assign g23 = 116'b00000000000000000000000000011111111111111111111111111111001111011111100000000000000000000000000000000000000000000000;
assign g24 = 116'b00000000000000000000000000011111111111111111111111111111011111011111111000000000000000000000000000000000000000000000;
assign g25 = 116'b00000000000000000000000000011111111111111111111111111111011110011111111111111111111111111000000000000000000000000000;
assign g26 = 116'b00000000000000000000000000011111111111111111111111111111011110111111111111111111111111111111111000000000000000000000;
assign g27 = 116'b00000000000000000000000000011111111111111111110000111111011110111111111111111111111111111111111111000000000000000000;
assign g28 = 116'b00000000000000000000000000011111111111111111100000011111011100111111111111111111111111111111111111110000000000000000;
assign g29 = 116'b00000000000000000000000000011111111111111111000000011111001101111111111111111111111111111111111111111100000000000000;
assign g30 = 116'b00000000000000000000111111101111111111111111000000011111000001111111111111111111111111111111111111111110000000000000;
assign g31 = 116'b00000000000000000001111111111111111111111111100000011111100011111111111111111111111111111111111111111111000000000000;
assign g32 = 116'b00000000000000000000111111111111111111111111111001111111111111111111111111111111111111111111111111111111100000000000;
assign g33 = 116'b00000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000;
assign g34 = 116'b00000000000000010000000000001111111111111111111111111111111111111111111111111111111111111110000000011111000000000000;
assign g35 = 116'b00000000000000111100000000001111111111111111111111111111111111111111111111111111111111111110000000000000000000000000;
assign g36 = 116'b00000000000000111100000000000111111111111111111111111111111111111111111111111111111111111111111111111110000000000000;
assign g37 = 116'b00000000000000111000000000000011111111100000000000000000000001111111111111111111111111111111111111111111111100000000;
assign g38 = 116'b00000000000001111000000000000001111100000001111111111000000011111111111111111111111111111111111111111111111111000000;
assign g39 = 116'b00000000000001111000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111100000;
assign g40 = 116'b00000000000000111000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111110000;
assign g41 = 116'b00000000000000110000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111110000;
assign g42 = 116'b00000000000000000001111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111110000;
assign g43 = 116'b00000000000000000011111100011111111100011111111100001111111111000111111111111111111111111111111111111111111111110000;
assign g44 = 116'b00000000000000000111111110001111111100011111111110000111111111000011111111111111111111111111111111111111111111100000;
assign g45 = 116'b00000000000000000001111110001111111110001111111111000111111111100011111111111111111111111111111111111111111111000000;
assign g46 = 116'b00000000000000000000000000000010011110001111111111100111111111110001111111111111111111111111111111111111110000000000;
assign g47 = 116'b11110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign g48 = 116'b11111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000111111111;
assign g49 = 116'b11111111111111111111111111111111111111111110000000000000000100011110010111100010000011100000111100001111111111111111;
assign g50 = 116'b11111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign g51 = 116'b11111111000111111111111111111111111100000011100111000111111111111111111111111111111111111111101111111111111111111111;
assign g52 = 116'b11111111000001111111100000001110000000000000000000000011111110011111001111111111111111111110000001111111100000000111;

always @(posedge clk) begin
    if(col > g_col && col <= g_col+116 && row > g_row && row <=g_row + 52)begin
		case(row-g_row)
        0 : nflag <= g1[116-(col-g_col)];
		1 : nflag <= g2[116-(col-g_col)];
		2 : nflag <= g3[116-(col-g_col)];
		3 : nflag <= g4[116-(col-g_col)];
		4 : nflag <= g5[116-(col-g_col)];
		5 : nflag <= g6[116-(col-g_col)];
		6 : nflag <= g7[116-(col-g_col)];
		7 : nflag <= g8[116-(col-g_col)];
		8 : nflag <= g9[116-(col-g_col)];
		9 : nflag <= g10[116-(col-g_col)];
		10 : nflag <= g11[116-(col-g_col)];
		11 : nflag <= g12[116-(col-g_col)];
		12 : nflag <= g13[116-(col-g_col)];
		13 : nflag <= g14[116-(col-g_col)];
		14 : nflag <= g15[116-(col-g_col)];
		15 : nflag <= g16[116-(col-g_col)];
		16 : nflag <= g17[116-(col-g_col)];
		17 : nflag <= g18[116-(col-g_col)];
		18 : nflag <= g19[116-(col-g_col)];
		19 : nflag <= g20[116-(col-g_col)];
		20 : nflag <= g21[116-(col-g_col)];
		21 : nflag <= g22[116-(col-g_col)];
		22 : nflag <= g23[116-(col-g_col)];
		23 : nflag <= g24[116-(col-g_col)];
		24 : nflag <= g25[116-(col-g_col)];
		25 : nflag <= g26[116-(col-g_col)];
		26 : nflag <= g27[116-(col-g_col)];
		27 : nflag <= g28[116-(col-g_col)];
		28 : nflag <= g29[116-(col-g_col)];
		29 : nflag <= g30[116-(col-g_col)];
		30 : nflag <= g31[116-(col-g_col)];
		31 : nflag <= g32[116-(col-g_col)];
		32 : nflag <= g33[116-(col-g_col)];
		33 : nflag <= g34[116-(col-g_col)];
		34 : nflag <= g35[116-(col-g_col)];
		35 : nflag <= g36[116-(col-g_col)];
		36 : nflag <= g37[116-(col-g_col)];
		37 : nflag <= g38[116-(col-g_col)];
		38 : nflag <= g39[116-(col-g_col)];
		39 : nflag <= g40[116-(col-g_col)];
		40 : nflag <= g41[116-(col-g_col)];
		41 : nflag <= g42[116-(col-g_col)];
		42 : nflag <= g43[116-(col-g_col)];
		43 : nflag <= g44[116-(col-g_col)];
		44 : nflag <= g45[116-(col-g_col)];
		45 : nflag <= g46[116-(col-g_col)];
		46 : nflag <= g47[116-(col-g_col)];
		47 : nflag <= g48[116-(col-g_col)];
		48 : nflag <= g49[116-(col-g_col)];
		49 : nflag <= g50[116-(col-g_col)];
		50 : nflag <= g51[116-(col-g_col)];
		51 : nflag <= g52[116-(col-g_col)];
        endcase
end
end

always@(posedge halfsec or posedge rst)begin
    if(rst) gflag<=0;
    else if(yb_flag == 1) gflag<=1;
    else gflag<=0;
end
//------------------------------------//fg
always@(posedge halfsec or posedge rst) begin
    if(rst) fg<=0;
    else if(yb_flag==2 && Flag && move == 1 && fg != 2) fg<=1; //��ܸ��D����}����
    else if(yb_flag==0 && fg && move == 1) fg<=2; //��ܸ��D�����F�ĤG�����D
	else if(move == 2) fg<=0;//���nn�����F
  //  else if(fg==2 && gg_row>=414 && move == 2) fg<=0;
    else fg<=fg;
end

//gg_row
always@(posedge halfsec or posedge rst) begin
	if(rst) begin
		gg_row<=414;
		move<=0;
	end
	else if(fg==2) begin
			if(gg_row>50 && (move == 0 || move == 1))begin
				gg_row<=gg_row-3;
				move<=1;
			end
			else if(gg_row<=50 && move == 1)begin
				gg_row<=gg_row;
				move<=2;
			end
			else if(gg_row<=50 && move == 2)begin
				gg_row<=gg_row+3;
				move<=move;
			end
			else if(gg_row>50 && gg_row<414 && move == 2)begin
				gg_row<=gg_row+3;
				move<=move;
			end
			else if(gg_row>=414 && move == 2)begin
				gg_row<=gg_row;
				move<=0;
				Flag<=0;
			end
			else gg_row<=gg_row;
	end
	else if(Flag == 1)begin
		 if(gg_row>174 && (move == 0 || move == 1))begin
				gg_row<=gg_row-3;
				move<=1;
			end
			else if(gg_row<=174 && move == 1)begin
				gg_row<=gg_row;
				move<=2;
			end
			else if(gg_row<=174 && move == 2)begin
				gg_row<=gg_row+3;
				move<=move;
			end
			else if(gg_row>174 && gg_row<414 && move == 2)begin
				gg_row<=gg_row+3;
				move<=move;
			end
			else if(gg_row>=414 && move == 2)begin
				gg_row<=gg_row;
				move<=0;
				Flag<=0;
			end
			else gg_row<=gg_row;
			
	end
		
	else if(yb_flag == 0) Flag<=1;
	else begin 
		gg_row<=gg_row; Flag<=Flag; 
	end
end

//////////////
wire [0:86*87-1] m_brick={
	87'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	87'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	87'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	87'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	87'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	87'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	87'b000000000000000000000000110000000000000000000000000000000000001000000000000000000000000,
	87'b000000000000000000000000111000000000000000000000000000000000011000000000000000000000000,
	87'b000000000000000000000000111100000000000000000000000000000000011000000000000000000000000,
	87'b000000000000000000000000111110000000000000000000000000000000111000000000000000000000000,
	87'b000000000000000000000000111111000000000000000000000000000001111000000000000000000000000,
	87'b000000000000000000000000111111110000000000000000000000000011111000000000000000000000000,
	87'b000000000000000000000000111111111000000000000000000000000111111000000000000000000000000,
	87'b000000000000000000000000111111111100000000000000000000011111111000000000000000000000000,
	87'b000000000000000000000000111111111110000000000000000000011111111100000000000000000000000,
	87'b000000000000000000000000111111111111100000000000000000111111111100000000000000000000000,
	87'b000000000000000000000001111111111111100000000000000001111111111100000000000000000000000,
	87'b000000000000000000000001111111111100000000000000000011111111111100000000000000000000000,
	87'b000000000000000000000001111111110000000000000000001111111111111100000000000000000000000,
	87'b000000000000000000000001111111100000001111111111001111111111111100000000000000000000000,
	87'b000000000000000000000001111110000011111111111111001111111111111100000000000000000000000,
	87'b000000000000000000000001111000011111111111111111101111111111111100000000000000000000000,
	87'b000000000000000000000001110000111111111111111111111111111111111100000000000000000000000,
	87'b000000000000000000000001100011111111111111111111111111111111111100000000000000000000000,
	87'b000000000000000000000000000111111111111111111111111111111111111100000000000000000000000,
	87'b000000000000000000000000001111111111111111111111111011111111111100000000000000000000000,
	87'b000000000000000000000000011111111111111111111111111110111111111000000000000000000000000,
	87'b000000000000000000000000111111111111111111111111111111101110000000000000000000000000000,
	87'b000000000000000000000001111111111111111111111111111111110000000000000000000000000000000,
	87'b000000000000000000000001111111111111111111111111111111111110001100000000000000000000000,
	87'b000000000000000000000011111111111111111111111111111111111111111110000000000000000000000,
	87'b000000000000000000000011111111111111111111111111111111111111111100000000000000000000000,
	87'b000000000000000000000111111111111111111111111111111111111111111001111000000000000000000,
	87'b000000000000000111000111111111111111111111111111111111111111111011111111100000000000000,
	87'b000000000011111111001111111111111111111111111111111111111111110111111111111110000000000,
	87'b000000001111111110001111111111111111111111111111111111111111111111111111111111111000000,
	87'b000000000111111110011111111111111111111111111111111111111111111111111111111111111110000,
	87'b000000000011111110011111111111111100111111001111111111111111111111111111111111111100000,
	87'b000000000001111110011111111111111100111111001111111111111111111111111111111111111000000,
	87'b000000000000111100011111111111111111111111101111111111111111011111111111111111100000000,
	87'b000000000000011100111111111111111111111111111111111111111111011111111111111111000000000,
	87'b000000000000001100111111111111111111111111111111111111111111011111111111111110000000000,
	87'b000000000000001000111111111111111111111111111111111111111111101111111111111100000000000,
	87'b000000000000000000111111111111111111111111111111111111111111101111111111111000000000000,
	87'b000000000000000000111111111111111111111111111111111111111111110111111111110000000000000,
	87'b000000000000000000111111111111111111111111111111111111111111110011111111100000000000000,
	87'b000000000000000000111111111111111111111111111111111111111111111000111111000000000000000,
	87'b000000000000000000111111111111111111111111111111111111111111111100000000000000000000000,
	87'b000000000000000000111111111111111111111111111111111111111111111110000000000000000000000,
	87'b000000000000000000111111111111111111111111111111111111111111111111110000000000000000000,
	87'b000000000000000000011111111111111111111111111111111111111111111111111000000000000000000,
	87'b000000000000000000011111111111111111111111111111111111111111111111111000000000000000000,
	87'b000000000000000000011111111111111111111111111111111111111111111111110000000000000000000,
	87'b000000000000000000001111111111111111111111111111111111111111111111110000000000000000000,
	87'b000000000000000000001111111111111111111111111111111111111111111111100000000000000000000,
	87'b000000000000000000000111111111111111111111111111111111111111111111100000000000000000000,
	87'b000000000000000000000111111111111111111111111111111111111111111111100000000000000000000,
	87'b000000000000000000000011111111111111111111111111111111111111111111111000000000000000000,
	87'b000000000000000000000011111111111111111111111111111111111111111111111110000000000000000,
	87'b000000000000000000000001111111111111111111111111111111111111111111111110000000000000000,
	87'b000000000000000000000000111111111111111111111111111111111111111111111111000000000000000,
	87'b000000000000000000000000011111111111111111111111111111111111111111111111100000000000000,
	87'b000000000000000000000000111111111111111111111111111111111111111111111111110000000000000,
	87'b000000000000000000000000111111111111111111111111111111111111111111111111110000000000000,
	87'b000000000000000000000001111111111111111111111111111111111111111111111111110000000000000,
	87'b000000000000000000000001111111111111111111111111111111111111111111111111100000000000000,
	87'b000000000000000000000001111111111111111111111111111111111111111111111111111000000000000,
	87'b000000000000000000000001111111111111111111111111111111111111111111111111111000000000000,
	87'b000000000000000000000011111111111111111111111111111111111111111111111111111000000000000,
	87'b000000000000000000000011111111111111111111111111111111111111111111111111100000000000000,
	87'b000000000000000000000011111111111111111111111111111111111111111111111111100000000000000,
	87'b000000000000000000000011111111111111111111111111111111111111111111111111111000000000000,
	87'b000000000000000000000011111111111111111111111111111111111111111111111111100000000000000,
	87'b000000000000000000000011111111111111111111111111111111111111111111111111111000000000000,
	87'b000000000000000000000011111111111111111111111111111111111111111111111111111000000000000,
	87'b000000000000000000000001111111111111111111111111111111111111111111111111111000000000000,
	87'b000000000000000000000001111111111111111111111111111111111111111111111111110000000000000,
	87'b000000000000000000000001111111111111111111111111111111111111111111111111100000000000000,
	87'b000000000000000000000000111111111111111111111111111111111111111111111111000000000000000,
	87'b000000000000000000000000011111111111111111111111111111111111111111111111000000000000000,
	87'b000000000000000000000000011111111111111111111111111111111111111111111100000000000000000,
	87'b000000000000000000000000001111111111111111111111111111111111111111110000000000000000000,
	87'b000000000000000000000000000111111111111111111111111111111111111111100000000000000000000,
	87'b000000000000000000000000000000111111111111111111111111111111111110000000000000000000000,
	87'b000000000000000000000000000000001111111111111111111111111111111000000000000000000000000,
	87'b000000000000000000000000000000000000000111111111111111111100000000000000000000000000000
};

assign brick = (m_brick[(row-414)*87+(col-bk_col)])? 1:0;
assign brick1 = (m_brick[(row-414)*87+(col-bk_col1)])? 1:0;
assign brick2 = (m_brick[(row-414)*87+(col-bk_col2)])? 1:0;
assign brick3 = (m_brick[(row-414)*87+(col-bk_col3)])? 1:0;
assign brick4 = (m_brick[(row-414)*87+(col-bk_col4)])? 1:0;

/////////////
//pixel_col
always@(posedge clk or posedge rst) begin 
	if(rst) pixel_col<=0;
	else if(pixel_col==H_pw) pixel_col<=0;
	else pixel_col<=pixel_col+1;
end

//pixel_row
always@(posedge clk or posedge rst) begin
	if(rst) pixel_row<=0;
	else if(pixel_col==H_pw) pixel_row<=pixel_row+1;
	else if(pixel_row==V_pw)pixel_row<=0;
	else pixel_row<=pixel_row;
end

//cnt
always@(posedge clk or posedge rst)begin
	if(rst) cnt <= 0;
	else if(cnt==25000000) cnt <= 0;//�b��
	else cnt <= cnt+1;
end

//counter
always@(posedge clk or posedge rst ) begin
	if(rst) counter<=0;
	else if(counter == 781250) counter<=0;
	else counter<=counter+1;
end

//random
always@(posedge clk or posedge rst ) begin
	if(rst) random<=0;
	else random<=random+1;
end


//day
always@(posedge clk or posedge rst ) begin
	if(rst) day<=SUN;
	else if(s_col<=0) day<=MOON;
	else if(m_col<=0) day<=SUN;
	else day<=day;
end
//s_col
always@(posedge clk or posedge rst ) begin
	if(rst) s_col<=400;
	else if(cnt == 781250 && day == SUN) s_col<=s_col-5;
	else if(s_col<=0) begin
		s_col<=800;
	end	
	else s_col<=s_col;
end
//m_col
always@(posedge clk or posedge rst ) begin
	if(rst) m_col<=800;
	else if(cnt == 781250 && day == MOON) m_col<=m_col-5;
	else if(m_col<=0) begin
		m_col<=800;
	end	
	else m_col<=m_col;
end
//up_col
always@(posedge clk or posedge rst ) begin
	if(rst) up_col<=800;
	else if(counter == 781250 && up_cho) up_col<=up_col-3;//�b���99pixel??
	else if(up_col<=0) up_col<=800;
	else up_col<=up_col;
end
//c_col
always@(posedge clk or posedge rst ) begin
	if(rst) c_col<=800;
	else if(counter == 781250 && c_cho && !invincible) c_col<=c_col-3;//�b���99pixel??
	else if(c_col<=0 || invincible) c_col<=800;
	else c_col<=c_col;
end

//bk_col
always@(posedge clk or posedge rst ) begin
	if(rst) bk_col<=799;
	else if(counter == 781250 && bk_cho[0]) bk_col<=bk_col-3;//�b���99pixel??
	//else if(counter == 781250 ) bk_col<=bk_col-3;//�b���99pixel??
	else if(bk_col<=0) bk_col<=799;
	else bk_col<=bk_col;
end

//bk_col1
always@(posedge clk or posedge rst ) begin
	if(rst) bk_col1<=799;
	else if(counter == 781250 && bk_cho[1]) bk_col1<=bk_col1-3;//�b���99pixel??
	else if(bk_col1<=0) bk_col1<=799;
	else bk_col1<=bk_col1;
end
//bk_col2
always@(posedge clk or posedge rst ) begin
	if(rst) bk_col2<=800;
	else if(counter == 781250 && bk_cho[2]) bk_col2<=bk_col2-3;//�b���99pixel??
	else if(bk_col2<=0) bk_col2<=800;
	else bk_col2<=bk_col2;
end
//bk_col3
always@(posedge clk or posedge rst ) begin
	if(rst) bk_col3<=800;
	else if(counter == 781250 && bk_cho[3]) bk_col3<=bk_col3-3;//�b���99pixel??
	else if(bk_col3<=0) bk_col3<=800;
	else bk_col3<=bk_col3;
end
//bk_col4
always@(posedge clk or posedge rst ) begin
	if(rst) bk_col4<=800;
	else if(counter == 781250 && bk_cho[4]) bk_col4<=bk_col4-3;//�b���99pixel??
	else if(bk_col4<=0) bk_col4<=800;
	else bk_col4<=bk_col4;
end
//timer
always@(posedge clk or posedge rst) begin
	if(rst) timer<=0;
	else if(choose && timer<5 && cnt == 25000000) timer <= timer+1;
	else if(timer == 5 ) timer<=0;//�ֿn���ӻ�ê��
	else timer<=timer;
end

//choose,choose2,bk_cho,up_cho
always@(posedge clk or posedge rst ) begin
	if(rst) begin
		choose<=0;
		choose2<=0;
		choose3<=0;
		bk_cho<=0;
		bk_num<=0;
		c_cho<=0;
		up_cho<=0;
	end	
	else if(cnt == 25000000) begin//�b��M�w�@��
		case(random)
			0,20,35:begin 
				choose<=1;
				bk_cho[timer]<=1;
			end
			45:begin
				choose3<=1;
				c_cho<=1;
			end	
			60:begin
				choose2<=1;
				up_cho<=1;
			end
			default:begin
				choose<=0;
				choose2<=0;
				choose3<=0;

			end	
		endcase
	end
	else if(bk_col<=0) begin
		bk_cho[0]<=0;
		bk_num<=bk_num+1;
	end
	else if(bk_col1<=0) begin
		bk_cho[1]<=0;
		bk_num<=bk_num+1;
	end	
	else if(bk_col2<=0) begin
		bk_cho[2]<=0;
		bk_num<=bk_num+1;
	end
	else if(bk_col3<=0) begin
		bk_cho[3]<=0;
		bk_num<=bk_num+1;
	end
	else if(bk_col4<=0) begin
		bk_cho[4]<=0;
	end
    else if(up_col<=0) begin
		up_cho<=0;
	end
	else if(invincible) c_cho<=0;
	else bk_cho<=bk_cho;
end

//gameover 
always@(posedge clk or posedge rst) begin
	if(rst) begin 
		gameover<=0; 
		life<=5; 
	end
	else if(!invincible) begin
		if(life == 0) gameover<=1;
		else if(col > gg_col && col <= gg_col+91 && row > gg_row && row <=gg_row + 87&& nnflag &&bk_cho[0] && brick & (col >= bk_col & col < bk_col+87 )&row>=414 & row<500 & row>=g_row & row<=g_row+52 & col>=g_col & col<=g_col+116 & nflag) life<=life-1;//����Ǫ�0
		else if(col > gg_col && col <= gg_col+91 && row > gg_row && row <=gg_row + 87&& nnflag &&bk_cho[1] && brick1 & (col >= bk_col1 & col < bk_col1+87 )&row>=414 & row<500 & row>=g_row & row<=g_row+52 & col>=g_col & col<=g_col+116 & nflag) life<=life-1;//����Ǫ�1
		else if(col > gg_col && col <= gg_col+91 && row > gg_row && row <=gg_row + 87&& nnflag &&bk_cho[2] && brick2 & (col >= bk_col2 & col < bk_col2+87 )&row>=414 & row<500 & row>=g_row & row<=g_row+52 & col>=g_col & col<=g_col+116 & nflag) life<=life-1;//����Ǫ�2
		else if(col > gg_col && col <= gg_col+91 && row > gg_row && row <=gg_row + 87&& nnflag &&bk_cho[3] && brick3 & (col >= bk_col3 & col < bk_col3+87 )&row>=414 & row<500 & row>=g_row & row<=g_row+52 & col>=g_col & col<=g_col+116 & nflag) life<=life-1;//����Ǫ�3
		else if(col > gg_col && col <= gg_col+91 && row > gg_row && row <=gg_row + 87&& nnflag &&bk_cho[4] && brick4 & (col >= bk_col4 & col < bk_col4+87 )&row>=414 & row<500 & row>=g_row & row<=g_row+52 & col>=g_col & col<=g_col+116 & nflag) life<=life-1;//����Ǫ�4
		else if(col > gg_col && col <= gg_col+91 && row > gg_row && row <=gg_row + 87&& nnflag &&row >= 400 & row < 430 & col >= up_col & col < up_col+100 & up_cho & row>=g_row & row<=g_row+52 & col>=g_col & col<=g_col+116 & nflag) life<=life-1; //upper brick
		else gameover<=gameover;
	end
	else gameover<=gameover;
end

//invincible,t_invincible
always@(posedge clk or posedge rst) begin
	if(rst) begin 
		invincible<=0;
		t_invincible<=0;
	end	
	else if(col > gg_col && col <= gg_col+91 && row > gg_row && row <=gg_row + 87&& nnflag && c_cho && candy &&row>= 320 & row < 400 & col >= c_col & col < c_col+84 ) invincible<=1;
	else if( invincible && cnt == 25000000 ) t_invincible<=t_invincible+1;
	else if( t_invincible==10 ) begin
		invincible<=0;
		t_invincible<=0;
	end
	else invincible<=invincible;
end
//row_a,row_b
always@(posedge clk or posedge rst) begin
	if(rst) begin
		row_a<=104'h5061737365643a303000;//Passed:00
		row_b<=104'h52656d61696e3a353000;//Remained:50
	end	
	//else row_a<=row_a;
	else begin
		row_a[43:40]<=quo;
		row_a[35:32]<=bk_bum-quo*10;
		row_b[43:40]<=quo1;
		row_b[35:32]<=20-(bk_bum-quo*10);
	end
end

//blink
always@(posedge clk or posedge rst)begin
	if(rst) blink<=0;
	else if(cnt == 25000000) blink<=~blink;
	else blink<=blink;
end

//color
always@(posedge clk) begin
	if(rst) color<=0;
	else if(visible) begin
		if (bk_num >= 20 && (!gameover)) color<=win;
		else if(gameover) color<=gg;
		//if((col-s_col)*(col-s_col)+(row-150)*(row-150)<=6400) color<=3'b110;//sun yellow 
        else if(col > gg_col && col <= gg_col+91 && row > gg_row && row <=gg_row + 87&& nnflag && !gflag)//body cyan
		begin
			if(invincible)begin
				if(blink) color<=3'b111;
				else color<=3'b100;
			end
			else color<=3'b100;
		end
        else if(col >= gg_col + 39 && col <= gg_col+61 && row >= gg_row+13 && row <= gg_row+20 && !nnflag && !gflag)color<=3'b110; // eyes
        else if(col >= gg_col + 45 && col <= gg_col+60 && row >= gg_row+31 && row <= gg_row+43 && !nnflag && !gflag)color<=3'b110;// buttons
        else if(col > g_col && col <= g_col+116 && row > g_row && row <=g_row + 52 && nflag && gflag) color<=3'b001;
		else if(row>= 270 & row < 350 & col >= c_col & col < c_col+84 & c_cho ) begin//candy
			if((row-c_row)>=25 & (row-c_row)<=46 & (col-c_col)>=22 & (col-c_col)<=59 & !candy) color<=3'b111;//���x red
			else if(candy) color<=3'b101;//face pink
			else begin
				case(day)
					SUN:color<=3'b011;//sky cyan
					MOON:color<=3'b001;//sky blue
			endcase
			end
		end 
		else if(row >= 100 & row < 300) begin//day
			case(day)
				SUN: begin
					if((col-s_col)*(col-s_col)+(row-200)*(row-200)<=10000) color<=3'b110;//sun yellow 
					else color<=3'b011;//sky cyan
				end
				MOON: begin
					if((col-m_col)*(col-m_col)+(row-200)*(row-200)<=10000) color<=3'b111;//moon white
					else color<=3'b001;//sky blue
				end
			endcase
		end
		else if(row >= 400 & row < 430 & col >= up_col & col < up_col+100 & up_cho)//upbrick white
		begin
			if(row>=405 & row<415 & col>=up_col+20 & col<up_col+50) color<=3'b000;
			else color<=3'b000;
		end
		
		//else if((row-310)*(row-310) +(col- c_col)*(col- c_col)<=81) color<=3'b101;//face pink
		else if(row>=414 & row<500 ) begin//bricks
			if(bk_cho[0] & (col >= bk_col & col < bk_col+87 )) begin
				if((row-414)>=37 & (row-414)<=39 & (col-bk_col)>=34 & (col-bk_col)<=43 & !brick ) color<=3'b000;//eyes black
				else if(brick) color<=3'b010;//green
				else color<=3'b110;
			end
			else if (bk_cho[1] & (col >= bk_col1 & col < bk_col1+87 )) begin
				if((row-414)>=37 & (row-414)<=39 & (col-bk_col1)>=34 & (col-bk_col1)<=43 & !brick1 ) color<=3'b000;//eyes black
				else if(brick1) color<=3'b111;//white
				else color<=3'b110;
			end
			else if (bk_cho[2] & (col >= bk_col2 & col < bk_col2+87 )) begin
				if((row-414)>=37 & (row-414)<=39 & (col-bk_col2)>=34 & (col-bk_col2)<=43 & !brick2 ) color<=3'b000;//eyes black
				else if(brick2) color<=3'b100;//red
				else color<=3'b110;
			end
			else if (bk_cho[3] & (col >= bk_col3 & col < bk_col3+87 )) begin
				if((row-414)>=37 & (row-414)<=39 & (col-bk_col3)>=34 & (col-bk_col3)<=43 & !brick3 ) color<=3'b000;//eyes black
				else if(brick3) color<=3'b001;//blue
				else color<=3'b110;
			end
			else if (bk_cho[4] & (col >= bk_col4 & col < bk_col4+87 )) begin
				if((row-414)>=37 & (row-414)<=39 & (col-bk_col4)>=34 & (col-bk_col4)<=43 & !brick4 ) color<=3'b000;//eyes black
				else if(brick4) color<=3'b101;//pink
				else color<=3'b110;
			end
			else color<=3'b110;
		end
		else if(row>= 500 & row < 600) color<=3'b000;//lower platform black 
		else if(row>= 0 & row < 400) begin
			case(day)
				SUN:color<=3'b011;//sky cyan
				MOON:color<=3'b001;//sky blue
			endcase
		end
		else if(row>= 400 & row < 600) color<=3'b110;//ground yellow
		else color<=3'b111;//white for debugging �]���z�פW�Τ���o��
	end
	else color<=3'b000;//black
end

endmodule
